library ieee;
use     ieee.std_logic_1164.all;

package GitVersionPkg is
   constant GIT_VERSION_C : std_logic_vector(31 downto 0) := x"34e82993";
end package GitVersionPkg;
